ENTITY device IS
	PORT(
		a, b: IN std_logic;
		y: OUT std_logic);
END device;