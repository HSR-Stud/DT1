LIBRARY library_name_1 {, libary_name_2; ...};
USE library_name.element_name;
--oder
USE library_name.ALL
--Beispiel
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;