signal identifier [, identifier, ...]: TYPE [:= value];
signal sig1, sig2: bit;
